`ifndef COMMON_VH
`define COMMON_VH
`define code_path "./code.txt"
`define data_path "./data.txt"
`define output_path "output.txt"

`define INIT_PC 32'h00003000
typedef logic [31:0] Vec32;
typedef logic [5:0] Vec6;
typedef logic [4:0] Vec5;
typedef logic [1:0] Vec2;
typedef logic [2:0] Vec3;
typedef logic [32:0] Vec33;
typedef logic [25:0] Vec26;
typedef logic [15:0] Vec16;

typedef enum Vec6 {
    ALU_ADD = 6'b100000,
    ALU_ADDU = 6'b100001,
    ALU_SUB = 6'b100010,
    ALU_SUBU = 6'b100011,
    ALU_LSHIFT = 6'b000000,
    ALU_LRSHIFT = 6'b000010,
    ALU_ARSHIFT = 6'b000011,
    ALU_LSHIFTV = 6'b000100,
    ALU_LRSHIFTV = 6'b000110,
    ALU_ARSHIFTV = 6'b000111,
    ALU_AND = 6'b100100,
    ALU_OR = 6'b100101,
    ALU_XOR = 6'b100110,
    ALU_NOR = 6'b100111,
    ALU_SLT = 6'b101010,
    ALU_SLTU = 6'b101011
} AluOp;

typedef enum Vec32 {
    ADD     = 32'b000000_????????????????????_100000,
    ADDU    = 32'b000000_????????????????????_100001,
    SUB     = 32'b000000_????????????????????_100010,
    SUBU    = 32'b000000_????????????????????_100011,
    SLL     = 32'b000000_????????????????????_000000,
    SRL     = 32'b000000_????????????????????_000010,
    SRA     = 32'b000000_????????????????????_000011,
    SLLV    = 32'b000000_????????????????????_000100,
    SRLV    = 32'b000000_????????????????????_000110,
    SRAV    = 32'b000000_????????????????????_000111,
    AND     = 32'b000000_????????????????????_100100,
    OR      = 32'b000000_????????????????????_100101,
    XOR     = 32'b000000_????????????????????_100110,
    NOR     = 32'b000000_????????????????????_100111,
    SLT     = 32'b000000_????????????????????_101010,
    SLTU    = 32'b000000_????????????????????_101011,

    ADDI    = 32'b001000_????????????????????_??????,
    ADDIU   = 32'b001001_????????????????????_??????,
    ANDI    = 32'b001100_????????????????????_??????,
    ORI     = 32'b001101_????????????????????_??????,
    XORI    = 32'b001110_????????????????????_??????,
    SLTI    = 32'b001010_????????????????????_??????,
    SLTIU   = 32'b001011_????????????????????_??????,

    LUI     = 32'b001111_????????????????????_??????,

    MULT    = 32'b000000_????????????????????_011000,
    MULTU   = 32'b000000_????????????????????_011001,
    DIV     = 32'b000000_????????????????????_011010,
    DIVU    = 32'b000000_????????????????????_011011,
    MFHI    = 32'b000000_????????????????????_010000,
    MTHI    = 32'b000000_????????????????????_010001,
    MFLO    = 32'b000000_????????????????????_010010,
    MTLO    = 32'b000000_????????????????????_010011,

    BEQ     = 32'b000100_????????????????????_??????,
    BNE     = 32'b000101_????????????????????_??????,
    BLEZ    = 32'b000110_????????????????????_??????,
    BGTZ    = 32'b000111_????????????????????_??????,
    BGEZ    = 32'b000001_?????00001??????????_??????,
    BLTZ    = 32'b000001_?????00000??????????_??????,

    JR      = 32'b000000_????????????????????_001000,
    JALR    = 32'b000000_????????????????????_001001,
    J       = 32'b000010_????????????????????_??????,
    JAL     = 32'b000011_????????????????????_??????,

    LB      = 32'b100000_????????????????????_??????,
    LBU     = 32'b100100_????????????????????_??????,
    LH      = 32'b100001_????????????????????_??????,
    LHU     = 32'b100101_????????????????????_??????,
    LW      = 32'b100011_????????????????????_??????,
    SB      = 32'b101000_????????????????????_??????,
    SH      = 32'b101001_????????????????????_??????,
    SW      = 32'b101011_????????????????????_??????,

    SYSCALL = 32'b000000_????????????????????_001100,
    NOP     = 32'b000000_00000000000000000000000000
} InstructionCode;

typedef struct packed {
    InstructionCode instructionCode;
    Vec5 rs, rt, rd;
    Vec16 imm16;
    Vec26 imm26;
    Vec6 funct;
    Vec5 shamt;
} Instruction;

typedef Vec5 GprID;

typedef enum Vec3{
    gprRegisterSrc_RS,
    gprRegisterSrc_RT,
    gprRegisterSrc_RD,
    gprRegisterSrc_RA, // 31
    gprRegisterSrc_R0  // 0
} GprRegisterSrc; // GprInput/WriteRegister

typedef enum Vec3{
    pipelineStage_IF_ID,
    pipelineStage_DECODE,
    pipelineStage_ID_EX,
    pipelineStage_EXECUTE,
    pipelineStage_EX_MEM,
    pipelineStage_MEMORY,
    pipelineStage_MEM_WB,
    pipelineStage_NEVER
}PipelineStage;

typedef enum Vec3{
    gprWriteInputSrc_imm16_lshift_16,   // valid in IF_ID_REG
    gprWriteInputSrc_pc_add_8,          // valid in ID_EX_REG
    gprWriteInputSrc_aluResult,         // valid in EX_DM_REG
    gprWriteInputSrc_mduResult,         // valid in EX_DM_REG
    gprWriteInputSrc_dmResult           // valid in DM_WB_REG
} GprWriteInputSrc;

function PipelineStage readyPipelineStage(GprWriteInputSrc gprWriteInputSrc);
    case(gprWriteInputSrc)
        gprWriteInputSrc_imm16_lshift_16: readyPipelineStage = pipelineStage_IF_ID;
        gprWriteInputSrc_pc_add_8: readyPipelineStage = pipelineStage_ID_EX;
        gprWriteInputSrc_aluResult: readyPipelineStage = pipelineStage_EX_MEM;
        gprWriteInputSrc_mduResult: readyPipelineStage = pipelineStage_EX_MEM;
        gprWriteInputSrc_dmResult: readyPipelineStage = pipelineStage_MEM_WB;
    endcase
endfunction

typedef enum Vec3{
    aluMduInputSrc_gpr1,
    aluMduInputSrc_gpr2,
    aluMduInputSrc_unsigned_imm16,
    aluMduInputSrc_signed_imm16,
    aluMduInputSrc_unsigned_shamt
} AluMduInputSrc;

typedef enum Vec2{
    // pcJumpMode_next, // jumpEnabled = 0
    pcJumpMode_rel, // beq
    pcJumpMode_abs, // j
    pcJumpMode_reg  // ja
}PcJumpMode;

typedef enum Vec2{
    // pcJumpInputSrc_pc_add_4,
    pcJumpInputSrc_gpr_read1,
    pcJumpInputSrc_signed_imm16_lshift_2,
    pcJumpInputSrc_unsigned_imm26_lshift_2
}PCJumpInputSrc;

typedef enum Vec3{
    pcJumpCondition_false,  // jumpEnabled = 0
    pcJumpCondition_true,
    pcJumpCondition_eq,
    pcJumpCondition_ne,
    pcJumpCondition_le,
    pcJumpCondition_lt,
    pcJumpCondition_gt,
    pcJumpCondition_ge
}PcJumpCondition;

typedef enum Vec3{
    dmReadType_unsigned_4 = 0,
    dmReadType_unsigned_1,
    dmReadType_signed_1,
    dmReadType_unsigned_2,
    dmReadType_signed_2
    // dmReadType_signed_4
}DmReadType;

typedef enum Vec2{
    dmWriteType_0, // no write
    dmWriteType_1,
    dmWriteType_2,
    dmWriteType_4
}DmWriteType;

typedef struct packed{
    GprRegisterSrc gprReadIDSrc1;
    GprRegisterSrc gprReadIDSrc2;
    PipelineStage gprResultRequiredStage1;
    PipelineStage gprResultRequiredStage2;
    GprRegisterSrc gprWriteIDSrc;
    logic gprWriteEnabled;
    GprWriteInputSrc gprWriteInputSrc;
    // PipelineStage gprWriteReadyStage; = dmWriteType == dmWriteType_0 ? 
    AluMduInputSrc aluMduInputSrc1;
    AluMduInputSrc aluMduInputSrc2;
    AluOp aluOp;
    // mdu related
    // dm always write from gpr read2
    DmReadType dmReadType;
    DmWriteType dmWriteType;
    PcJumpMode pcJumpMode;
    PCJumpInputSrc pcJumpInputSrc;
    PcJumpCondition pcJumpCondition;
}ControlSignal;

`define getGprID(RESULT, GPR_REGISTER_SRC, INSTRUCTION) \
    case(GPR_REGISTER_SRC) \
        gprRegisterSrc_RS: RESULT = INSTRUCTION.rs; \
        gprRegisterSrc_RT: RESULT = INSTRUCTION.rt; \
        gprRegisterSrc_RD: RESULT = INSTRUCTION.rd; \
        gprRegisterSrc_RA: RESULT = 5'b11111; \
        gprRegisterSrc_R0: RESULT = 5'b00000; \
    endcase

`define init_instruction(INSTRUCTION) \
    INSTRUCTION.instructionCode = NOP; \
    INSTRUCTION.rs = 5'b00000; \
    INSTRUCTION.rt = 5'b00000; \
    INSTRUCTION.rd = 5'b00000; \
    INSTRUCTION.imm16 = 16'b0000000000000000; \
    INSTRUCTION.imm26 = 26'b00000000000000000000000000; \
    INSTRUCTION.funct = 6'b000000; \
    INSTRUCTION.shamt = 5'b00000;

`define init_instruction_unblocking(INSTRUCTION) \
    INSTRUCTION.instructionCode <= NOP; \
    INSTRUCTION.rs <= 5'b00000; \
    INSTRUCTION.rt <= 5'b00000; \
    INSTRUCTION.rd <= 5'b00000; \
    INSTRUCTION.imm16 <= 16'b0000000000000000; \
    INSTRUCTION.imm26 <= 26'b00000000000000000000000000; \
    INSTRUCTION.funct <= 6'b000000; \
    INSTRUCTION.shamt <= 5'b00000;

`define init_control_signal(CONTROL_SIGNAL) \
    CONTROL_SIGNAL.gprReadIDSrc1 = gprRegisterSrc_R0; \
    CONTROL_SIGNAL.gprReadIDSrc2 = gprRegisterSrc_R0; \
    CONTROL_SIGNAL.gprResultRequiredStage1 = pipelineStage_NEVER; \
    CONTROL_SIGNAL.gprResultRequiredStage2 = pipelineStage_NEVER; \
    CONTROL_SIGNAL.gprWriteIDSrc = gprRegisterSrc_R0; \
    CONTROL_SIGNAL.gprWriteEnabled = 1'b0; \
    CONTROL_SIGNAL.gprWriteInputSrc = gprWriteInputSrc_aluResult; \
    CONTROL_SIGNAL.aluMduInputSrc1 = aluMduInputSrc_gpr1; \
    CONTROL_SIGNAL.aluMduInputSrc2 = aluMduInputSrc_gpr2; \
    CONTROL_SIGNAL.aluOp = ALU_ADD; \
    CONTROL_SIGNAL.dmReadType = dmReadType_unsigned_4; \
    CONTROL_SIGNAL.dmWriteType = dmWriteType_0; \
    CONTROL_SIGNAL.pcJumpMode = 'bx; \
    CONTROL_SIGNAL.pcJumpInputSrc = 'bx; \
    CONTROL_SIGNAL.pcJumpCondition = pcJumpCondition_false;

`define init_control_signal_unblocking(CONTROL_SIGNAL) \
    CONTROL_SIGNAL.gprReadIDSrc1 <= gprRegisterSrc_R0; \
    CONTROL_SIGNAL.gprReadIDSrc2 <= gprRegisterSrc_R0; \
    CONTROL_SIGNAL.gprResultRequiredStage1 <= pipelineStage_NEVER; \
    CONTROL_SIGNAL.gprResultRequiredStage2 <= pipelineStage_NEVER; \
    CONTROL_SIGNAL.gprWriteIDSrc <= gprRegisterSrc_R0; \
    CONTROL_SIGNAL.gprWriteEnabled <= 1'b0; \
    CONTROL_SIGNAL.gprWriteInputSrc <= gprWriteInputSrc_aluResult; \
    CONTROL_SIGNAL.aluMduInputSrc1 <= aluMduInputSrc_gpr1; \
    CONTROL_SIGNAL.aluMduInputSrc2 <= aluMduInputSrc_gpr2; \
    CONTROL_SIGNAL.aluOp <= ALU_ADD; \
    CONTROL_SIGNAL.dmReadType <= dmReadType_unsigned_4; \
    CONTROL_SIGNAL.dmWriteType <= dmWriteType_0; \
    CONTROL_SIGNAL.pcJumpMode <= 'bx; \
    CONTROL_SIGNAL.pcJumpInputSrc <= 'bx; \
    CONTROL_SIGNAL.pcJumpCondition <= pcJumpCondition_false;


typedef struct packed {
    Vec32 pcValue;
    Instruction instruction;
} IF_ID_REG; 

typedef struct packed {
    Vec32 pcValue;
    Instruction instruction;
    ControlSignal controlSignal;
    Vec5 gprReadRegister1;
    Vec5 gprReadRegister2;
    Vec5 gprWriteRegister;
    Vec32 gprWriteInput;
    Vec32 gprResult1;
    Vec32 gprResult2;
} ID_EX_REG;

typedef struct packed {
    Vec32 pcValue;
    Instruction instruction;
    ControlSignal controlSignal;
    Vec5 gprReadRegister1;
    Vec5 gprReadRegister2;
    Vec5 gprWriteRegister;
    Vec32 gprWriteInput;
    Vec32 gprResult1;
    Vec32 gprResult2;
    Vec32 aluResult;
    Vec32 memoryForwardingResult1;
    Vec32 memoryForwardingResult2;
    logic memoryForwardingEnabled1;
    logic memoryForwardingEnabled2;
} EX_MEM_REG;


typedef struct packed {
    Vec32 pcValue;
    Instruction instruction;
    ControlSignal controlSignal;
    Vec5 gprReadRegister1;
    Vec5 gprReadRegister2;
    Vec5 gprWriteRegister;
    Vec32 gprWriteInput;
    Vec32 gprResult1;
    Vec32 gprResult2;
    Vec32 dmReadResult;
} MEM_WB_REG;

`endif